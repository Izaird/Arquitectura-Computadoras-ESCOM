----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:25:13 02/27/2019 
-- Design Name: 
-- Module Name:    Sumador1 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Sumador1 is
    Port ( a,b,cin : in  STD_LOGIC;
           suma,cout : out  STD_LOGIC);
end Sumador1;

architecture Behavioral of Sumador1 is
begin
	suma<=a xor b xor cin;
	cout<= (a and b) or (b and cin) or (a and cin);
end Behavioral;

